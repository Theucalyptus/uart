../clkUnit/clkUnit.vhd